module circuit(
    input A,
    output B
);

assign B = ~A;

endmodule